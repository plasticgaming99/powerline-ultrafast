module main

import os

const colorrune_cap_small = 16
const colorrune_cap_mid = 48
const colorrune_cap_large = 192

fn colorify(s string, cfg string, cbg string) []ColorRune {
    mut cr := []ColorRune{cap: colorrune_cap_small}
    for r in s.runes() {
        cr << ColorRune{
            fg: cfg
            bg: cbg
            text: r
        }
    }
    return cr
}

fn (mut cr1 []ColorRune) joincrs(cr2 []ColorRune) {
    if cr1.len == 0 {
        cr1 = cr2.clone()
        return
    }
    mut fg := ""
    if cr1.last().bg != "1" {
        fg = cr1.last().bg
    } else {
        fg = cr2.first().bg
    }
    joint := colorify(pl_symbol, fg, cr2.first().bg)
    cr1 << joint
    cr1 << cr2
}

fn (mut cr1 []ColorRune) joincrs_right(cr2 []ColorRune) {
    mut cr := []ColorRune{cap: colorrune_cap_mid}
    if cr1.len == 0 {
        cr1 = cr2.clone()
        return
    }
    if cr2.len == 0 {
        return
    }
    joint := colorify(pl_symbol_r, cr1.last().bg, cr2.first().bg)
    //cr1.insert(0,joint)
    //cr1.insert(0, cr2)
    cr << cr2
    cr << joint
    cr << cr1
    cr1 = cr.clone()
}

fn (mut cr1 []ColorRune) draw_right(cr2 []ColorRune) {
    mut i2 := 0
    for i := cr1.len - cr2.len; i < cr1.len; i++ {
        cr1[i] = cr2[i2]
        i2++
    }
}

fn (mut cr []ColorRune) add_padding(val int) {
    mut p := cr[0]
    p.text = ` `
    mut f := cr.last()
    f.text = ` `
    cr.insert(0, p)
    cr << f
}

struct Username{
}

fn (username &Username) getrunes() []ColorRune {
    mut cr := []ColorRune{cap: colorrune_cap_small}
    lname := os.loginname() or {"unknown"}
    cr = colorify(lname, user_fg, user_bg)
    cr.add_padding(padding)
    return cr
}

struct Hostname{
}

fn (hostname &Hostname) getrunes() []ColorRune {
	mut cr := []ColorRune{cap: colorrune_cap_small}
    cr = colorify(os.hostname() or {"unknown"}, host_fg, host_bg)
    cr.add_padding(padding)
    return cr
}

struct Cwd {
}

//fn (cr []ColorRune) joindircr([]ColorRune) {

//}

fn (cwd &Cwd) getrunes() []ColorRune {
    mut cr := []ColorRune{cap: colorrune_cap_mid}
    mut inhome := false
    mut inroot := false
    mut rootstr := "/"
    //mut dirtrunc := 0
	wd := os.getwd()
    hd := os.home_dir()
    ws := wd.split(os.path_separator)[1..]
    hs := hd.split(os.path_separator)[1..]
    if ws.len > 1 {
        if ws[hs.len-1] == hs[hs.len-1] {
            inhome = true
        }
    }
    $if windows {
        if wd.runes()[1] == `:` {
            inroot = true
            rootstr = wd.runes()[..2].string()
        }
    } $else {
        if wd == "/" {
            inroot = true
        }
    }


    if inhome {
       mut c := colorify("~", home_fg, home_bg)
       c.add_padding(padding)
       cr << c
       if ws.len == hs.len {
        return cr
       }
    } else if inroot {
       if ws[0] == "" {
          mut c := colorify(rootstr, path_fg, path_bg)
          c.add_padding(padding)
          cr << c
          return cr
       }
    }

    mut cr2 := []ColorRune{}

    if inhome {
        for i, s in ws[hs.len..] {
            mut c := []ColorRune{}
            if i == ws.len-hs.len-1 {
                c = colorify(s, cwd_fg, path_bg)
            } else {
                c = colorify(s, path_fg, path_bg)
            }

            c.add_padding(padding)
            if i != 0 {
                mut c2 := colorify(separator, path_fg, path_bg)
                cr2 << c2
            }
            cr2 << c
        }
        cr.joincrs(cr2)
    } else {
        for i, s in ws {
            mut c := []ColorRune{}
            if i == ws.len-1 {
                c = colorify(s, cwd_fg, path_bg)
            } else {
                c = colorify(s, path_fg, path_bg)
            }

            c.add_padding(padding)
            if i != 0 {
                mut c2 := colorify(separator, path_fg, path_bg)
                cr2 << c2
            }
            cr2 << c
        }
        cr.joincrs(cr2)
    }

    return cr
}

// end dollar or percentage $ %
struct PromptEnd {
}

fn (pe &PromptEnd) getrunes() []ColorRune {
    mut cr := []ColorRune{cap: colorrune_cap_small}
	cr << ColorRune{
        bg: cmd_passed_bg,
        fg: cmd_passed_fg,
        text: prompt_end.runes().first(),
    }
    cr.add_padding(1)
    return cr
}

